#Initial commit
#Store main code here
